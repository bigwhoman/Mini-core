module CU(
input [1:0] op,
input clk,


output halted,
output data_mem_write
);



endmodule